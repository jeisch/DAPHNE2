-- endpoint.vhd
-- master clock distribution for DAPHNE2 includes Bristol Timing Endpoint Logic
-- 
-- MMCM0: takes 100MHz system clock and produces SCLK100, SCLK200, local 62.5MHz clock
--        this MMCM is reset by a hard reset from the uC
--
-- MMCM1: choose between local 62.5MHz clock or timing endpoint 62.5MHz clock. Generates the master clock 62.5MHz
--        and fast clock 437.5MHz for the front end. use_ep is the bit that does the switching.
--
-- Timestamp is generated by endpoint (use_ep=1) or faked with free running counter (use_ep=0)

-- jamieson olsen <jamieson@fnal.gov>

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity endpoint is
port(

    sysclk_p, sysclk_n: in std_logic; -- system clock LVDS 100MHz from local oscillator
    reset_async: in std_logic; -- async hard reset from the microcontroller

    -- external optical timing SFP link interface

    cdr_sfp_los: in std_logic; -- loss of signal
    cdr_sfp_abs: in std_logic; -- high if module is absent
    cdr_sfp_tx_dis: out std_logic; -- high to disable timing SFP TX
    cdr_sfp_tx_p, cdr_sfp_tx_n: out std_logic; -- send data upstream (optional)

    -- external CDR chip interface

    adn2814_clk_p, adn2814_clk_n: in std_logic; -- LVDS recovered clock 312.5MHz
    adn2814_data_p, adn2814_data_n: in std_logic; -- LVDS recovered serial data 
    adn2814_los: in std_logic; -- loss of signal
    adn2814_lol: in std_logic; -- loss of lock

    -- timing endpoint interface 

    ep_reset: in std_logic; -- soft reset endpoint logic
    ep_edgesel: in std_logic; -- sample CDR data on rising or falling edge of CDR clock
    ep_addr: in std_logic_vector(7 downto 0); -- Endpoint address (async, sampled in clk domain)
	ep_tgrp: in std_logic_vector(1 downto 0); -- Timing group (async, sampled in clk domain)
    ep_ts_rdy: out std_logic; -- endpoint timestamp is good
    ep_stat: out std_logic_vector(3 downto 0); -- endpoint state bits

    -- misc interface signals

    mmcm1_reset: in std_logic;
    mmcm1_locked: out std_logic;
    mmcm0_locked: out std_logic;

    use_ep: in std_logic; -- 0 = run on local clocks with fake timestamp, 1 = use endpoint clocks and real timestamp

    mclk: out std_logic;  -- master clock 62.5MHz
    fclk: out std_logic;  -- fast clock for frontend
    sclk200: out std_logic; -- system clock 200MHz
    sclk100: out std_logic; -- system clock 100MHz

    timestamp: out std_logic_vector(63 downto 0) -- sync to mclk

  );
end endpoint;

architecture endpoint_arch of endpoint is

component pdts_endpoint_stdlogic
port(
		sclk: in std_logic; -- Free-running system clock
		srst: in std_logic; -- System reset (sclk domain)
		addr: in std_logic_vector(7 downto 0); -- Endpoint address (async, sampled in clk domain)
		tgrp: in std_logic_vector(1 downto 0); -- Timing group (async, sampled in clk domain)
		stat: out std_logic_vector(3 downto 0); -- Status output (sclk domain)
		rec_clk: in std_logic; -- CDR recovered clock from timing link
		rec_d: in std_logic; -- CDR recovered data from timing link (rec_clk domain)
		sfp_los: in std_logic := '0'; -- SFP LOS line (async, sampled in sclk domain)
		cdr_los: in std_logic := '0'; -- CDR LOS line (async, sampled in sclk domain)
		cdr_lol: in std_logic := '0'; -- CDR LOL line (async, --sampled in sclk domain)
        pll_locked: in std_logic;
		clk: out std_logic; -- 50MHz clock output
		rst: out std_logic; -- 50MHz domain reset
		rdy: out std_logic; -- Timestamp valid flag
		sync: out std_logic_vector(3 downto 0); -- Sync command output (clk domain)
		sync_stb: out std_logic; -- Sync command strobe (clk domain)
		sync_first: out std_logic; -- Sync command valid flag (clk domain)
		tstamp: out std_logic_vector(63 downto 0); -- Timestamp out
		debug: out std_logic_vector(31 downto 0); -- port for debug info, e.g. applied delay values
		txd: out std_logic;
		tx_dis: out std_logic);
end component;

signal sysclk_ibuf: std_logic;
signal mmcm0_clkfbout, mmcm0_clkfbout_buf: std_logic;
signal mmcm0_clkout0, mmcm0_clkout1, mmcm0_clkout2: std_logic;
signal local_clk62p5: std_logic;
signal sclk100_i: std_logic;

signal adn2814_clk_ibuf, adn2814_clk: std_logic;
signal adn2814_data: std_logic;
signal ep_rec_d_ddr: std_logic_vector(1 downto 0);
signal ep_rec_d: std_logic;

signal ep_clk62p5: std_logic;
signal cdr_sfp_txd: std_logic;

signal mmcm1_clkfbout, mmcm1_clkfbout_buf: std_logic;
signal mmcm1_clkout0, mmcm1_clkout1, mmcm1_clkout2: std_logic;
signal mclk_i: std_logic;

signal real_timestamp, fake_timestamp, timestamp_reg: std_logic_vector(63 downto 0);

begin

-- sysclk is 100MHz LVDS, receive it with IBUFDS. sysclk comes in on bank 33
-- which has VCCO=1.5V. IOSTANDARD is LVDS and the termination resistor is external (DIFF_TERM=FALSE)

sysclk_ibufds_inst : IBUFGDS port map(O => sysclk_ibuf, I => sysclk_p, IB => sysclk_n);

mmcm0_inst: MMCME2_ADV
generic map(
    BANDWIDTH            => "OPTIMIZED",
    CLKOUT4_CASCADE      => FALSE,
    COMPENSATION         => "ZHOLD",
    STARTUP_WAIT         => FALSE,
    DIVCLK_DIVIDE        => 1,
    CLKFBOUT_MULT_F      => 10.000, -- VCO = 1000MHz
    CLKFBOUT_PHASE       => 0.000,
    CLKFBOUT_USE_FINE_PS => FALSE,
    CLKOUT0_DIVIDE_F     => 16.000, -- CLKOUT0 = 62.5MHz
    CLKOUT0_PHASE        => 0.000,
    CLKOUT0_DUTY_CYCLE   => 0.500,
    CLKOUT0_USE_FINE_PS  => FALSE,
    CLKOUT1_DIVIDE       => 5, -- CLKOUT1 = 200MHz
    CLKOUT1_PHASE        => 0.000,
    CLKOUT1_DUTY_CYCLE   => 0.500,
    CLKOUT1_USE_FINE_PS  => FALSE,
    CLKOUT2_DIVIDE       => 10, -- CLKOUT2 = 100MHz
    CLKOUT2_PHASE        => 0.000,
    CLKOUT2_DUTY_CYCLE   => 0.500,
    CLKOUT2_USE_FINE_PS  => FALSE,
    CLKIN1_PERIOD        => 10.000 -- 100MHz system clock input
)
port map(
    CLKFBOUT            => mmcm0_clkfbout,
    CLKFBOUTB           => open,
    CLKOUT0             => mmcm0_clkout0, -- 62.5MHz
    CLKOUT0B            => open,
    CLKOUT1             => mmcm0_clkout1, -- 200MHz
    CLKOUT1B            => open,
    CLKOUT2             => mmcm0_clkout2, -- 100MHz
    CLKOUT2B            => open,     
    CLKOUT3             => open, 
    CLKOUT3B            => open,
    CLKOUT4             => open,
    CLKOUT5             => open,
    CLKOUT6             => open,
    CLKFBIN             => mmcm0_clkfbout_buf,
    CLKIN1              => sysclk_ibuf,
    CLKIN2              => '0',
    CLKINSEL            => '1', -- high to use CLKIN1
    DADDR               => (others=>'0'),
    DCLK                => '0',
    DEN                 => '0',
    DI                  => (others=>'0'),
    DO                  => open,
    DRDY                => open,
    DWE                 => '0',
    PSCLK               => '0',
    PSEN                => '0',
    PSINCDEC            => '0',
    PSDONE              => open,
    LOCKED              => mmcm0_locked,
    CLKINSTOPPED        => open,
    CLKFBSTOPPED        => open,
    PWRDWN              => '0',
    RST                 => reset_async
);

mmcm0_clkfb_inst: BUFG port map( I => mmcm0_clkfbout, O => mmcm0_clkfbout_buf);

mmcm0_clk0_inst:  BUFG port map( I => mmcm0_clkout0, O => local_clk62p5); -- local clock 62.5MHz

mmcm0_clk1_inst:  BUFG port map( I => mmcm0_clkout1, O => sclk200); -- system clock 200MHz

mmcm_clk2_inst:  BUFG port map( I => mmcm0_clkout2, O => sclk100_i);  -- system clock 100MHz

sclk100 <= sclk100_i;

-- 312 MHz recovered clock from ADN2814 chip

cdr_clk_ibuf_inst: IBUFDS
generic map( DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS_25" )
port map( I => adn2814_clk_p, IB => adn2814_clk_n, O  => adn2814_clk_ibuf );

cdr_clk_bufg_inst: BUFG
port map( I => adn2814_clk_ibuf, O => adn2814_clk );

-- serial recovered data from ADN2814 chip

cdr_data_inst: IBUFDS
generic map( DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS_25" )
port map( I => adn2814_data_p, IB => adn2814_data_n, O  => adn2814_data );

-- choose rising or falling edge of the 312.5MHz CDR clock to sample the CDR data....

-- Verilog from Adrian:
--    IDDR #(.DDR_CLK_EDGE ("SAME_EDGE_PIPELINED")) iddr_timing
--    (
--        .Q1 (ep_rec_d_ddr[0]),
--        .Q2 (ep_rec_d_ddr[1]),
--        .C  (adn2814_clk),
--        .CE (1'b1),
--        .D  (adn2814_data),
--        .R  (1'b0)
--    );   

IDDR_inst: IDDR
generic map(DDR_CLK_EDGE => "SAME_EDGE_PIPELINED", INIT_Q1 => '0', INIT_Q2 => '0', SRTYPE => "ASYNC")
port map(
    Q1 => ep_rec_d_ddr(0),
    Q2 => ep_rec_d_ddr(1),
    C => adn2814_clk,
    CE => '1',
    D => adn2814_data,
    R => '0',
    S => '0'
);

-- Verilog from Adrian:
-- always @(posedge adn2814_clk) ep_rec_d = ep_rec_d_ddr [edge_sel];

edge_sel_proc: process(adn2814_clk)
begin
    if rising_edge(adn2814_clk) then
        if (ep_edgesel='1') then
            ep_rec_d <= ep_rec_d_ddr(1);
        else
            ep_rec_d <= ep_rec_d_ddr(0);            
        end if;
    end if;
end process edge_sel_proc;

-- Bristol UK timing endpoint, legacy timing interface using 8b10b encoded stream @ 312.5Mbps

pdts_endpoint_inst: pdts_endpoint_stdlogic
port map(
    sclk => sclk100_i, -- 100MHz from MMCM0
	srst => ep_reset,
	addr => ep_addr,
	tgrp => ep_tgrp,
	stat => ep_stat,
	rec_clk => adn2814_clk,
	rec_d => ep_rec_d,
	sfp_los => cdr_sfp_los,
    cdr_los => adn2814_los,
	cdr_lol => adn2814_lol,
    pll_locked => '1', -- originally intended for external PLL, not used
	clk => ep_clk62p5, -- output clock from endpoint 62.5MHz
	rst => open, -- endpoint reset output not used here
	rdy => ep_ts_rdy,
	sync => open, -- sync commands not used by DAPHNE
	sync_stb => open,
	sync_first => open,
	tstamp => real_timestamp, -- this is sync to ep_clk62p5
	debug => open,
	txd => cdr_sfp_txd, 
	tx_dis => open
);

-- you can TRY to send endpoint data upstream....

OBUFDS_inst: OBUFDS
generic map(IOSTANDARD=>"LVDS_25")
port map( I => cdr_sfp_txd, O => cdr_sfp_tx_p, OB => cdr_sfp_tx_n );

-- ...but the timing SFP transmitter is DISABLED, so nope.

cdr_sfp_tx_dis <= '1';

-- MMCM1 chooses between local clock 62.5MHz or the endpoint clock 62.5MHz
-- after switching be sure to reset this MMCM! From the selected clock generate
-- the master 62.5MHz and the 437.5MHz clock needed for the front end

mmcm1_inst: MMCME2_ADV
generic map(
    BANDWIDTH            => "OPTIMIZED",
    CLKOUT4_CASCADE      => FALSE,
    COMPENSATION         => "ZHOLD",
    STARTUP_WAIT         => FALSE,
    DIVCLK_DIVIDE        => 1,
    CLKFBOUT_MULT_F      => 14.000, -- VCO = 875MHz
    CLKFBOUT_PHASE       => 0.000,
    CLKFBOUT_USE_FINE_PS => FALSE,
    CLKOUT0_DIVIDE_F     => 2.000, -- CLKOUT0 = 437.5MHz
    CLKOUT0_PHASE        => 0.000,
    CLKOUT0_DUTY_CYCLE   => 0.500,
    CLKOUT0_USE_FINE_PS  => FALSE,
    CLKOUT1_DIVIDE       => 14, -- CLKOUT1 = 62.5MHz
    CLKOUT1_PHASE        => 0.000,
    CLKOUT1_DUTY_CYCLE   => 0.500,
    CLKOUT1_USE_FINE_PS  => FALSE,
    CLKOUT2_DIVIDE       => 14,
    CLKOUT2_PHASE        => 0.000,
    CLKOUT2_DUTY_CYCLE   => 0.500,
    CLKOUT2_USE_FINE_PS  => FALSE,
    CLKIN1_PERIOD        => 16.000 -- CLKIN1 = 62.5MHz 
)
port map(
    CLKFBOUT            => mmcm1_clkfbout,
    CLKFBOUTB           => open,
    CLKOUT0             => mmcm1_clkout0,  -- 437.5MHz
    CLKOUT0B            => open,
    CLKOUT1             => mmcm1_clkout1,  -- 62.5MHz
    CLKOUT1B            => open,
    CLKOUT2             => open, 
    CLKOUT2B            => open,     
    CLKOUT3             => open, 
    CLKOUT3B            => open,
    CLKOUT4             => open,
    CLKOUT5             => open,
    CLKOUT6             => open,
    CLKFBIN             => mmcm1_clkfbout_buf,
    CLKIN1              => ep_clk62p5,     -- endpoint clock 62.5
    CLKIN2              => local_clk62p5,  -- local clock 62.5
    CLKINSEL            => use_ep,         -- 1 = CLKIN1 = endpoint clock, 0 = CLKIN2 = local clock
    DADDR               => (others=>'0'),
    DCLK                => '0',
    DEN                 => '0',
    DI                  => (others=>'0'),
    DO                  => open,
    DRDY                => open,
    DWE                 => '0',
    PSCLK               => '0',
    PSEN                => '0',
    PSINCDEC            => '0',
    PSDONE              => open,
    LOCKED              => mmcm1_locked,
    CLKINSTOPPED        => open,
    CLKFBSTOPPED        => open,
    PWRDWN              => '0',
    RST                 => mmcm1_reset
);

mmcm1_clkfb_inst: BUFG port map( I => mmcm1_clkfbout, O => mmcm1_clkfbout_buf);

mmcm1_clk0_inst:  BUFG port map( I => mmcm1_clkout0, O => fclk); -- fast clock 437.5MHz for front end logic

mmcm1_clk1_inst:  BUFG port map( I => mmcm1_clkout1, O => mclk_i); -- master clock 62.5MHz

mclk <= mclk_i;

-- make a fake timestamp for when we're running with local clocks (use_ep=0) free running counter

fake_ts_proc: process(mclk_i)
begin
    if rising_edge(mclk_i) then
        if (reset_async='1') then
            fake_timestamp <= (others=>'0');
        else
            fake_timestamp <= std_logic_vector(unsigned(fake_timestamp) + 1);
        end if;
    end if;
end process fake_ts_proc;

-- mux and register the timestamps in the master clock domain
--
-- CDC WARNING! real_timestamp launches in ep_clk62p5 domain, but is captured in mclk domain.
-- IF the endpoint clock is selected (use_ep=1) THEN mclk and ep_clk62p5 are frequency locked.
-- BUT the phase is unknown due to routing delays and latency through MMCM1. It is possible 
-- that timestamp_reg may capture garbage here. We'll have to see and maybe make this CDC more robust...

ts_proc: process(mclk_i)
begin
    if rising_edge(mclk_i) then
        if (use_ep='1') then
            timestamp_reg <= real_timestamp; -- from endpoint
        else
            timestamp_reg <= fake_timestamp;
        end if;
    end if;
end process ts_proc;

timestamp <= timestamp_reg;

end endpoint_arch;
